//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
N1OpbXnm5z3qjRznMOym0a3GaQBkDvBiQUmV3+D8wPs5493IP5+oMt+MpTZPDTPs
TjLEILGY/H6Z574Y1r7qXP/15cTE0T+lLN5lYyz+EtLRSsl0qgGEz26jutB29ZST
y9UHYLNMoGCSW3j/vJPriQ3WbfsMLryB7aTcz3MVi+pIGLX3sljIKOugNOwmt6C2
dlq7tZ5jQOYrcG8k5VtGYZUzlmB19kOlHnn0OMP1LE+kmsYJt5JqZdOxbL+scZYF
qUCdYZWs+53H6XYwBMjlcoeFALnOJYsORV6oMF02w1y7zBopC2vjWwGyeOPIq0MS
fq/LNLHPfQA+4oTcYLGV5w==
//pragma protect end_key_block
//pragma protect digest_block
55LgwGH1AKY+lXBDwW+zTOz3RQQ=
//pragma protect end_digest_block
//pragma protect data_block
ho85RNpPuAfILX/4VLQariAPX+cKO48iX+U6FMq7jGRgzQ0RI0BOfRwuGioqH9JZ
70hff02wETBRESWl2UIOGO4/1iDmVAIr6AA8iW/n97NA5s+dA8hzkGpwvn0CSjRa
9DjmYUpaBBqq0RGkaYv27kSYHd022fQdd/8pndYnQUxCi/n2sLelgGJqV6/m2F2S
dEnWiZiAoaPh/fNgSvwDzcig9DehNmWRJmM3CzaSBENcPXDcv3e4QzyR8AUMyULd
Q9v60g4fGT4D4fKZ8TmTNoNMrDZmvuxEHJDAFc+MkY588GXYEB4kzSKGnFVb/l5H
zcyu9POqLpYselz2CpyBhh1XGkBNeSEC4fUCO3Bqk8G59wV+rNrFzK3XRHfhZly/
47HJm62j+DSRDAFOmI7MSF6fSJiNpQugF5RlLkHOhJ0uwfemfkhSj0cD0PCF6HVV
LIbXyUJ0UyyoLu3288ILCtFQ3oWrxANontr9ZItQ8C7c+r1UX3mtnQr1tIE1mcP4
J7rALFo4O63cFwnkSOp4Dlq34kwE9/sKoh9k7Wt4IiHoLzCIbj5ls6AXM0QZW2bI
JX+kgAMXhnB+FWvloTTnlKusWn7LGRgSrXfIHAegNcTVjg/vC340RzK2gUMGa+P3
cqlMlda5fG2ZZqWyCE59QfbeOfelSZnbv7CC6/6MOPT+ZNJbZ3HHPjpgZnOPcGZn
dX/9KurHBpk5TFm64Xsue2MpyR7fqdt6XLwT4AuP4s9bpl7ck+ME96nQ1EfbV77D
jjzw/EMjXzMCTMQUJXvEgEMxTYRiI4o/AhJZFw9bH0lC/UPyyGN5VW7cK2GPzefs
arV7jL4KrqNgb7xr5GJzg5TTmwLbRJg/rkc0ahPSQe5lekq0wY+41C9lBEH4wmgL
Q6ZdeH3ELHn889uv+AX4ODtB4CGstdthXBUbuHOpjM5jognqHCYeujxxuFCznMYC
gKQqwlyixsBepGknUcByWE/UwcavBpkKDbYwK/X0GURCUwG3bdHtXjOV4z37o1Tw
TWOASR9woHqH7+NVZtWgyhbtlb5WJUCcPjCId1Sh3PBkIL+af2FV/TaIUREfJOou
pjtK5EPyUdWzHOwLmaprQViCQyj/osD2WSsw5XnckJWuLqsUaVmZooJeZqdVDG7i
BEIIVXHGmnvj3s6U0wvXH8D5/bhS8ABTU094j4xaIOdDu0tQNpJIJjR6bEwzG5Bq
O8bfk5sTm34yoUSzq0rfnXEBOe8sygbl38NOKvNPa9V1re2vbX+2SldagfMVStiv
YS71/UQrfezBRCL3EOs8z5eRpAOgko+6bkNMaHLCEr1qYwVj7iVUdw+9C9DFoJjT
XpPNYfMsJd4z+e3/DKUi6ZNskaKGpKenRBo3rFwxCZT47hTsDalnALjmonhYQ0SZ
nL8vdMqoMKEjV9DSS+O4Hbh4DaCBBX6YXvFVx+UG6W3oDkfn9R3oXEmlpJUPf30t
P/yZnBxOgM1tsyXTDGyvkxhI/7a+mw/F5bOQ0/hSYmN8JfUsSrtQiNtOnzIAXGXk
yrD8XSWVm8yP9hRh729ZRE2rQz4isMsJP5GDCkIBU6prF/rOW0CnvK0PatpyP2+8
/Pv+3vBfcn5abjKUZnz8MaOstgFBQB6hryLDiANctxXoeHwLVJIMfuX0o0vGue0f
nTp48BGW4Ax1BtRIHfJHU6B2zCmXXMayenXfP6zmXGXa+5KEoczzoBDtiT8KspT7
I+rn9Vmrx9akK2hyBuKfAuuK1LXd7d+3q5Grx+3oVc65dtn1fXflQBltfBXAnPuS
KD15O+iKpTOvEt+NVq3Olf95zzuf6jZ9oyaUZeEmUx/6ivMwx4ICG4sxIu9ag9yj
1rWNAfZpXkZK5NbTO7AzplRdUxGdCuKZPvH4XYU/80sGr+207TnKimcgB87uWJMb
B/Z41/R2Lw77CtEtxU3dmsdB5Av/DIkmE/pcQnD5G6Ge63lmpRXLL9Uny3/2/YpG
D6LVkFDGixgbk4qFjrCllSYHnEnJSnkirn6tUd8P+X2Bc3YbKEjv5HZPNEVilD2c
xg0OBq3PLE5toeDjvGurWuMgEnVk69w/KLEmtkc1RVirxJmWUR1062QHTYWVwNJQ
YF+7VoWv/OxQj61RRsPi4Ty/mhCMI5ZpU9NhcuUBkvmSiDztqebk5ORXRadNnLrT
he6fgUttBwe7w4WsQiY6L8A0+TYS8Lp6mmtSmbJ++tazbvjPWXGL0Py+0Ipq4Hew
R4RnMJW+yTUYjcspJ4yUy6boOmb77DzxJHzHb1Odz37KaoEhsnGgdCE1kyxpOHPg
MWeR4UxM84+/cRWlBIQAPzyZWf2auqbI2rn8bYo93KxvLoWSUz93MAurjTBERPbj
5/bZ522brUOUyhurVimx6aDmxKS+Hdv8t9Kb88lQLiUTjSSjSRkAZWElBwXl55gX
Ut/1aeW0d4Mc23pjhEpwa9qQI8Lv8X19noH9dwFd/bpI5OW76z9rX3e6i2mmgwjs
BgilFwi0EY3kJaANGMJwk2jxF75AJPp9QD8SKFa30Yl+EZQNl1ESpaoLz7oykS5q
R15WpLVNbf4F1DTj9cmj6Bi6if76TAsJGwdFkfRT3rHt460PnKrI8/vWbnlv+z53
dyqXqQ6/NG0QxvJyECbNbAH9FagcGQp7KkIHaFSMVsYE4u8kSjpAK1LRgNjORJJa
uF6KEXnUzvnJc78ggGNQyzogj7RykLOnzLMOj7I6ztNxU3nJLSNFDbJvjExo8AP3
tnbo4oNFLeRLtoHFcUbiyPY81j+XqRRT15gICds3lIx1lX2mSbgeGNv4VWHjWpZq
qzOBWLMNKqI4AqZz83mGKuV/xtFf/faLwvKKKUhRkeB86xwr6MZ8cngFnEM7SFBq
OvlaRWUY2lwVsfnpq9JdfGDz6wxQoBVrbtbhUy8iL4rjARUi7dtQ730BTsQ9gq9C
WOuHMYuhP+zO9IXEBqiXv9Lq9RvfOJ2OgrGrdUz6LX1l5fO7Ias9msrcyN9fJQ8r
AQVaH+JQCr6lZ8dFlyu6nJJyx3JDztOsqQnNej1wCnUPGsSBcY6JSCohYa+Savpp
+uiybGg5ivzfG61USOd1eWkXYtv4h+WjPfDSBVObB2rhxhaRXvreh3/ShuhHhzYu
xD0C4N+IUlnO/AFekEvm2JY+jwLbdpJLL/ohSOOabLW1DeC/9NgWWOB96p/YOM0c
BFNbNIZYRXMomKp/h4DWRq49LkA+iNfW4D7cCn7TZKfjw4J5I3rwEbyi3dwTs+Vw
OTPlm25ermVVdGZIYh218GKSpyXv3a7M2hb38QfCdW3++P2jBBK2TKIXD+v87n4i
WeJFdOkSEi7RCAbeYzLXPS85buyJ/d7B9Q2A6+mea8gXTLLUlDLhqLVKmgyCxj6b
5P9sVsr6ZJAF2gMyBTr/Phv8KBQlv0Xk4FB3eR/AioH01mp1FT4AL7afaxpGVINR
lWiLEB7LKMyMOWDR57FiVByi+y961UfNc5CQeQIaFPvVcFF9vlMJkUPn1EMJ/E4U
+wbJlpOxzp8FHqxLphHrAulc09WVSQX/MIrAa+wxswSXoRaeO0OetfzJjh1X/MvI
vLIHXym/kTaM3iuO7YDcIP9pnQcsTRiA4Y3/Z8FrnJjy+7bxDPaSI+GbAH8ZIhlj
GbEX2c5pQsyfTQI2ke2W3Zip5D6DjvbhNf8xUFRG193lLrkXSx3dcinM5J/cRKUh
L4GNRE4hFg7H1i0c99WuGMrIco/jGB73T+94U2J4r/f8y4CgaAP1c6R3CQ3vbnk3
g/fDXil1auSQvWEW1mNDb7CytLzCxNqvrGsjtGFQl1lIONCrSCJpX3km7LydLwPU
q55rOS9eqvxIyKjWcbaw54ZUJHD8nhhbXqzVMrC2++hiL1FmYVlu+vn+5CYkIuef
zc2O0Ua2QzMnwiEeFbduUOL5Ee7w3RfMDEcEgBqXqjJ34Hmxwg53L/vRmDKd4Od7
dqh1gPo29O76sLQYHwty4BdEsGcTNi++F/qpdowoDwm3UTvnW2kdFDYr7So8hGuZ
CjYBAXuU/K0jQxfuTeHTZ0XmRZEe1aUfQ18A8D9BMp/8FyuJHICoDSvz2lf3qK5M
K9Al7JecVPXv68alrtNewFod3Lov+MLkK0r9W0qCoBWOrth+Q2yqIl8tCrswF4wo
2c7dTfJWlpYGZMt2p8W/trvLQ4Re4Zn6bFdwLTtXOxisnKpuTd7USnXrDc+0Cpbj
YTslKqo0QS2BYzhN7T7DkT1NOydAScBIYimSfTiDak+PpoQRzg7TtHN1E0qHOIuA
gYTRr9DywyN9wpJNzCLPh3Uygtncbbaz+1Mm7Eqtzc+aBiz9HfscsIdDH2ERH+rk
uf+MR1d/KrA3Qx685NYgqLY44qTEFYhJFUrcWpD3dxUKu8M5onolRAn9VLDZRHoE
CFRwMqE71suEA5dK4emlP4TZ1eRZVn8s4zdFzBPejWrV1ZvuQvETKDPT1YnGceJd
JS0fRsx7bR0pgGC+YiVvisRFM2U0gC3dUFt//zA9cdUcxmYJeYwALidTM5bkbiTd
Vq0XWKqH4VQqP8V48DU6x2wDyRk9UXriPyaqV60l3bcZe7iL7l1RvDAvA0MIeLFH
3fl++/wKE79eiQD+fuGqzRNw2uS7xgzkfyFXM7tZIsqUtSoypTeyzIn4yflBhRTl
c904SRHpHzA72uN4qqJb428rEcrXg9kf51UWxWeK0Ycjwp6DLMqZrQCvKslc6NH8
DBb6zifzQBnZ+RnZqkyTYYkfCxYgNQwzOs1TkXwf48kIE/VjH/8jHxccK9iorkFp
LbRVnhusnJjcT3D25OriS5JoYkJ8McaFTP9N+uqiI98nhlBVFAbmOIoJtqla1MRQ
oefIerhpgdKVYW+D0ZYMjk6GOQjp1kkCqXOz0+uWmLSBm8IQ7Q4pvJGxB9X+TIfs
ykPmHM2iroz0FraO9PYZKS9UkSapOw7yUVn3IAt0Pl91I37lnlNvlYf9/VSuOIeM
z9isCIEJP8PpYR+Qsei14DHGNFqFmryIz+uqrQR6jllWNdjlDDnga/7mdoLlV/o6
sC1HGLnQSTW54eAUvQfiJGiJiG/YvzatK4O0uTDoDtAVdaLMZDAgun1zmFPqB/8l
vYrmtLbz7jV2LxsX6D2LtOTr7bVa4dNTkKWmB+9wfWFZBgVA2C6YVNdrMZ9LMEfp
eX8ngIZOJZgEWTGVik0oWiodctwqaEgQzc2EGFF9qj+753WsoG54FYhsM7O30zcx
a4o4dsfLkBUetBZcn4PpToDqoC+3soggCT6iesixXuxnA7lxQkGkZHJ5DnvlHYHj
DYJ08zuwbVGoroVfiyK4wJe4s4R1YDxC8Zck/1gcAeXyeZIyo1foFUQMOM3X5Dj1
qxuMcyy0afM7lGD+17sS7Ap0wG0/WWk1uanzEWvip6ifWYiuqgXc1Ir6ku6NW8Hj
NNceCll9Gvb7J5oEWTV8OGUD/XSLYKp1e+qLJf/H0oykntfNT2ZXISHWltHOi0W0
a8hG+SawEdzRoCjS7J4PX/Tmj2b2icYUionRYeh4HBhL2lLnN3IgBojI9nZy+Lp7
7A3urFnlrHc3AOBblpOM5QbIhTnFSGVPwS/GWM9UFe5AlCxBcmZfV2zp1m2MQkV4
zRaPdzJDjMnKOmL2IKEp4d0limECi4W4CLs36dPjSjZh8QcabU0TcXUMmkkF6Mcz
+Qh2s3t1kOqA7SdxQ6aNnIBjWv30efwwwhzj3eoPqXYwxLlUac8vkrSIHiCSk8uf
J3yclW8GBGzOzCqUisoo+ZdCv8q6J1Jwrfr/XWn0lJpGUUtLC5XhslcGBFgMo58J
fm0ArvgUgX+hb768OE5xEOWbdCtDNqa3jGyhLzBoQGrdyiw1YL2eG3XXyudlEqFP
pw06jUjt+FTlsviy9dTbp6kB3bgjfEzY2Lwq8PjfltO9sRlno9N6BQ1duI/zy67p
IO130PGOM4h7qKZQj0kM6l0zF4QZUtn723Fte54Ez8+sC3Jq7Yub7rdWchc/8Oas
DalCD2m72EvGMGVIaUuk6EO81qjzJAZ4+pfZzrfFKlg6iLwb2EIlMBk4PgdAi2ou
8vNZR8xTq5WjH8E7pCcZ+YvJAj7q9CGGsZsg0zP5zRkn4D2JejZtzl9cWn8Au8wd
efGn/Mbq+ynmJsM2GpJIYBrvdDKyHXpNWsE7TpbghhFHnbvjPGy/h3J8tT+jhkqE
+iYSmderbW/FGQjDiuvA07jTon1Yg5I37Lpmy4f3Is+XCETBcfOv0dkvUbZwQ+0V
OVJFodNnJU1xHsEZy53QSkousEfEQdvXPEdo4DneGA5jXWvB7URc6jsBWa0Qbghi
Sl41ps6WUfqFKtL0JpuE9iYNjijlCghHnF8lJdw/r6fBCudPlwZis3l761FFClDj
bHk7Xf2g4lWCb9SI2PxJDakJsvH3E1KZmYs02xFQ8IBH+i7xOywfh9XTnhnP5EOl
NwGGmIwVa0+zkQzlh/4f9PFqVlZpDzHCxqu3Uf/DrPM1ET7S93UHHCcLyrNMEvg9
TPJ1yVmfgcewaQ0CdV5JXNc5ZKZA20V+Twc2KPKSKaRuzk9NgMH/WmczHjVYkmvw
6eo1HQSPH0iywd3GXk2fW/hnbUfU84ts0Xg1E2GJlE0CMIBjfFxoQpkA8GEraK+2
O+oaxtiMn+QaZ0JQaXnvb/9ZlTA+/AxGA2u9gDq8w+oHmAFq5ENOePEs0j6YN8wJ
1dSJxFGdfyLfkoMvASo5hgGxjvbCOwHyrokgAWAapGzsSDM2G4NGi5tggSw+dWDy
Fg5xCn22QVoB49F8fg2Jzc9L7mus/pQguGLqjRPozHjsoC8rnEsstWCM3zpib0bj
idOyOgnkTt+bWXMPWiDMFYkr6o37HbSOfE1dkZGFcMgyAkK0tUVPlnqWJrCLDV+E
iMOxQafno6IjjVfT2n87Jk/mkmZEXZgnyg1d/Bcg3zYKQaTZKfAUf5IlvhEcVmrL
KeDb0vdCHH8rarZxpUfdEpEoOb9xgO0PSUR68ixYDIc04ZCrvV9h7+gzYNQvPEnQ
/1Wiq/ZgoglbOtEdjqVmH1V+k8qjsXXlyUteO/cUq/+hMdUnhyqIAsp1/e6fSFMd
55RLt6VjDJ8VMrF75ONI0+NazO/c8bo8BEf5R9UoDJ7Z7V4+H79WfVWAAbKpqIv8
P7s2j7UkGsW9u3+2cbP3MBv1KDtT6BV0aREvTNqiNYAYd/shJv66c4Qx5zTc50xE
nCrDTp8GcNSC7pK4TS4YjQZOqeQCJQHGJVqnfLI5SCyTwN6+wk8I0UP+yyIID05t
kI/axGNeGdi2TNebQYFr9ilacY5Zwr+xvQco8luunGsfeD55SkrL972xM+2/2aNu
HZZaPhKn5DElkiHG0v6UEhPMUw+Nt6dlAMijVWM7JB7x3oh79hyHomcc6h6+Kw9m
Oq8lFAy39/YvP9JFyQ959aW71qjLLmG6czJT/8iUa6wzZiRk75KqQhwb4pYcRZ2C
e32WKpfEysnLbjY+yZoRCxPTKFg1bvQ1l5g/6J6H8st73IoVgO/9JbOwtX14Szlm
pPYOROy0XvPriMVfiWZ98xTsw5eZ1OnRHsZQu2FPDLeClQnd18e1iul9780R7nqX
OpXYGmxFlOLSJwwuL9GqR15CYiLhKHsgsP4M2gAEzJp5WYniKJtWk4AwALd2cmYl
xHtRrms9skd4OcXv5YVgDsdYxNbaXIomX6UqiB6mFm29YaWOjQAb5Xnq5MArH8+c
bIG8ASrus5ecElwQvp2EqW0g9QNV/b/2CXI+Ng5/gacRNM79l5ECWvaI9m978ceH
TQbwxKXxBWbKhyJpPzXbcTJAjJWYGaJwrHs2hHeg8uZwp9hMYmejDkf+oFkCe1Gs
7MzKi30EPd2zbMHkxAN084CwkY/r/VplLIrdTfOv3fEjzYlnIsdcuI4B1nEvDuyF
knAGZc0CjnQd6BraD8bMaaPOdi8t8/E7uO9Zz2z0Sk9lC2kjWTFxZ1nc8JeD60LB
LrwA99Wf48ci8xh/XkO4uOJTC3N2d0wZypkhq43JUHuAQ7rtQBd1m0DxEOXk/IiY
CTwLWLDB6N6pC4vs2onoYvwTb1b/SOd26g3vO3cIFF5QWG8/Uv6GbCAFSEjzzVzx
MUy9+KvHxnuAQn4z757upkBb5T2Wj8nHEyXbTeCGfxJ+p5rdUyB0VugDgWQyqxe8
G+PutkbMb28c1WiDpB1yj/PlWl4rfN9/nsY2DgxIXG+yDaZBoiRRPVrJxijzFJ8D
wr8/X7kRdwzjQaOl/UQ92kuC0Y1fvw+vCmivK+leecWN4YgPsI4AePvnD6jgkjHY
eeUN95C+c7oiT7c5fcHbXz0GjhWmz1xrnCYQKGkrKfwtvj+Qga+3ED2j0OCDj3Ua
wAqIVfwqNsQU5YbVOp0qDkVvsYpE0v5ieNFbMKJKwoWHQREOnyr3Ba7L+WtqOnO2
s9s4IKW9ittkP7z94bnfeyNfs11CSNX53uAxf2kKf7/TBAM9wXBDLJtEQ7D+54Uh
7gAXBfPMT6anHZLNK2DR0Rl3kAuGC/4XfWyyF6dta+qguKVkkgRK4q/DNtKCdIM/
yR3/nQybpuSE1obv8+LQGjFKZ+D+xzFB8DhxdtHneZvcM2uakmc/PorGhiJGfZ+K
9Gp8xYxHAlm/TEddua6Pqq8bIR+XLWMn/UDF8yjCeJK0SjUhhgf5p/iofnbbRw9+
gFXc65fI5K9IicSI7RE+CnBhcdtK5GO7UpyPFGosxJcdVH86+8+9NoUomVhAb2aO
Z8QCGuGLMHFRC5c13RiHXwj5oZrxU/azv33kkJQkvFx9rDMJasUS8tQD8QhQMiQv
EAYEVSxaRID9bmze6Yp3iUSapodO4fSFEeTqPTuBhIgFvlOgGLDm2yWx99emyHAP
P3SXpq3JubHUIGLBWV2PQIVmFDTfi7YqbNLlgxTSN+nTstVJm+RonlSwacxTQrCk
MEEkv75vDz0lyht1NwU8KBFX7o3Y61NErAicCFQuEZVrd6hz0LXu0oh3vkIWyhuY
C/wYfb0yBrZYUzt7d4mzCcxxwgeZ64lWSmzAjTIi/qrVD57E9BhCDvLE1iJqQDyW
+Z6uyUrcyeG/vDUskYuiJROZj3KuFHDk1LP+zGzudV2psoKqFfmQge/jsbcByw6l
QuwdX/7vWZHmtgS7znuT2hSviX6iz+hplnyM7k9CTyla7ZyBGLPWmlQxQhFbH3NA
vm6rybtNR4n9qxQdeD659lFl3W0UKE/+/cnNF1SAMC4W/nfLOx362TQyznuBklVV
NyhMCF9MjCOrFW3vCh7TJ+kp4BQH1LZbA5XW+uVdUJN+/fMYfBAQ21g714Ad1kui
RLF0tKWLwHwLmMiibVL7h29Bet/19ZeLi5DcR6xnclTgru69DojYX2ZlvTqLaiQQ
JWQNI/8U3NEOFFnpO6LFItUF7TyodibQ3djF+Mx+xoNfDw7YkkaGc6l9mALRBtJN
iZ0NhlWI3YAUfu9MS7JxfkGP5guSALENUFfFvZB0BlUAd+JAvxi2Bx4tbHZh/h3g
u0Lfxbk3Sgl2GTsv00QmKyXcAany1FdhkyONfo4vlFKp23ONvSg1auSkbOgikqX8
PRxhxds2leT+qKqr/5oP9h5l4u5E394hXcd20tuSRybbcpt37nWVCDW4s1zGIvLr
4/CReTsL9cgfYUF2ay8tvZEH3RdCpDuSCPczaEQQ0vt1zNU6u8l7wkmeuK+bP7V0
aO918Hv75AvxQ1L6wDQRoCUQu47hk6I6F7kNQOCOmTeXHJE/ux1jcK5XMUHOLUEp
uoRLLy8SOYtHhIhdqxxZfB9MlOxTSD9TV5I6LjHVYHsAK3DrkqFbnMvVQ9wNVUjG
LzqwcFI0dbkDF2LZW6p3RruS8mhNdLPcl+Kd5jOgcVMdSZPHU6gjfy+vbeiPrwkQ
rnBmAILRI7HyTunM91s145FqcOtBccoDoQ9/oeisaujVZ16CN3VM75pJwiuLooi/
PJg14xhg8iC89XDhi6V9MiIHxmRWfhN28Ern2ok3U0Lhe9NbUoIXUQkTTlBi5V2/
ei95DP0bzoNERAsAP29f0E9thAmjWEaATeVUQkb6ryiNJIGeD+UWqk/RhIcIpS6K
VrV1ypYUdk+F561UK/e9c1h8oww/RE35zfBhOl6sosUqgCTqsEtKm5v0zjrXIUML
x5F/1yc6tgUa/JFvIvbLAydMx7A3Q9oBgoKh2xwHqOSMhmDKk5/KlnfAHWnazEuU
3VKqCrqDQlgEF6axo3lohL8d5NOeRtDMhwJuG6C+dPj3s+Vh73eH/P85ZTmvna33
BTQuq6FMFt9BfIobXKRWJpzHueGcuZk0BweLm3IwPCA9Bio6MlYWdWSG4yw4fwYK
2ISk5yvKiJCm6SqaIREBDEwFgVpcbpcnee1UaGJPamhICgVL3rdm99JEdsOCHy4X
FzBtdMu1mfzrpROliasuUT26lRBUttQtqSt4EreB2hi8zkNJpbG+qpDuw96FBgzS
/glXdCXMFA5MPooYmPtRhnMKqVFIXGya/4SVQa13MfXR/CZ9+D/v3sLxvGvD1PhP
XTY0qVlGx1iU//xCaYZC86zhLsp4yyhfEloPxJURlkMs2BM6SYSlTNrqno4Xd0wJ
4+7p/4W0YyblIhnCitl+wNS6f05hWugQPkC8skhcLF8hAvYmla9v1hx2sS040F7v
9uQUdVmRgV2E7xMjuT5t+w2bBzW09ntAey0AJEFnqGrvIIsJLcEwTwvrMQpaspKy
bn2UcKT+uK8u0ukWVC4bvhmkJeajiv8lJC2Eqzp0qw6zAgbVC5UIMf22j7YtKZZ+
wy1ubPrn+H5iwqIzHml7YzCpE6mfmZDd6njX7djpfK91FSwLF1r8QhqbJ8PugWLp
5WcZspFK9E0WZ56RmcABRhJY5ihb/wMvVNYZ01OK9ATPYQeFbBkCUjedwo/k0gtb
TMH6CLUyK5QOUM5N5qxDqNwdmKwHgXHYhO836lcSISePScizBxzFIMs94wxTgSoE
FDT5b9K+1cdavv1pMF28b0aZtq0+a4rosb8c6qkRqKLAywiO6Uc38+Zkd5TEEkuj
VXVEcZ7GN3vKn/Z+v5yOdK9N6Wve2YcwNOUooyZmDZLSx0AiNWcmrLeT4lDHCK+f
RaqLmFnS3wuJb1YjKnjg7TpoC8hD5ZJxpn0W14pnrEbvospfCNyp8hr72jeL/bVH
s4SzLHKwglSdCxZYQumVbM4M6AEUm2Y6VmLyCiaoHQwpjV08qDGjvuWPh8Wte7RR
b1xea4Btc1c7EfPAaqLMPfprdNKnxlzqO8jvQpiIrylgQ/hl5CQtFet21waF6qAG
hKq9OJTCXn/q7A4ifTnjZYLzdvYyxYrNI61fCdzl53idQ9GgVr13FAcZreySb/cW
XZFEpqL5zH11Gtv+7MyhcExt35pH4I/RDE3jU88xaUtwvJ5EfFoMIeZMpPSsxeBW
cxL0PMd3u/wflyI6O6mE7vn7Ah1dU/EM5SCCFC0HS8jkcDRBzpqasR+eT+3jGYEb
D0Iz1I2RDvGYnKsVjX8mHwjh6ErayQWGljr8EHu6VQvE5CqmTgOPgSf+bDoLDQlm
xiofotab5bM7ICG5w/jt8GPsqMfIupWNL5CoURQtf4Sq8ZTtRM4PLfCfqVNu0o2M
tquE9Mgyo/B0BKay73PWftd3Vp2RHf1Kr37LFJy4lnrvZT69R46ayhnZP/lPUf+x
KE0SjGlEFEL53n6WLqRWc4MP/5UidTzWMX80INW7IEymj9s+LqM8MOKzDgal/LoA
y79QeJnQwGgP+/t66Yy6/jMxqJNlnOrsaeSliS0RfqEw+WmJeKrC+J0EBmTdbY1k
Cwf514EQeKNE/tHYiWqnqx63+Pgpws9lSHcIF4qioNlp6CNIbrSoVJWsNJ44dSVa
coJ0oSNA+FjJIkYs5A+o0EiD8oOc64rIb4hGMusDdx/IAOfObMW9s83wdm5xKFQw
jLoygQKeVqOeLAg8mGId+CUiByHKjxPQpR59wd1MU9uQgI18YB3k6cLAGhaxZifL
iOPMBUEXWYpi80Z3trvr3isyHLLqwekrPkvEn/Ekvs/+rbUpzraK8m7XB17/SJsw
XFS9qlaYhiX2wADOU3QM/JkQJrW9CeEIBNQaSlHyyClOEzDkESMpX/p7g7sVSmid
+LWIJ8SJJGBtpy0NnTdafoLkPhCDlBIWmSzZZhmGgiHQ/Gke7CMplKnO7aDbo15+
7m+CRWNufG7GAQrNwIqFKT/tw+oR8N/XsbGLwj8NmYnu42WrOI/+u9tl2F5Pjtrz
5t381nq++CCkwJriTUmHCYQbkEIZc4tVZs0nLlXnAdwZRByhMVFIwSWEbnL1tPWc
AcCIuYLS/4erKxq/6w7+neb3GlGnGOEXb8giYTOWqf5oZVn6RPZ+qi+TDp+i9P7G
cBI7Ej49z1yP+CyWAUeQe+sQN1+VqoohQkB+cfEBc4QDaC07fMYeGcl5mZK8LAXv
Z0Tphgz/qpkIvoZtlnfE2o7YpH00Robo5i2DWInF5Gbt+HQNyiJ9h9xmX5Rhf3XW
eGcrv+o3S/gMrPW4Uv72iwxDUrN4gw+dfHFjRKY0LzZKoqmOItAi7BqNSUyeM/4E
w/dBt2UEMjJkxghB3n/ne5gvpY0Y+P7xKenhHk0GlVGPfVxA0uWSWhCY4jGf0Zm9
/yzsSDOxa6/DNydvZFgDor4Hc80vMWf+4kpqbSJclGO79vKs/8LOOyEAV4dZZJZp
F0YZJJq/YjausxSQ76Bf8p+tGOf9/PhjQK7GxOTus2rJ39xifo2SzUMCfZrF/H/g
U0c4KykiRfDtiCLXfereCPuD0CPO7mMbzX3Kzcs1bRsdw+EbKA0SpxWTLimeOLW0
3oq2eL9yOUNWIKIfGgx3SRe6aTWfs0+VoDsXG1MoEd5fPuwB2SSlgiMx6Ly3WxtO
gKYOn7Vt2aMlA11ozBv0M8afMrenmOq5YpR/MOacQqx9mujj4WbTCTbjvUixHSvj
CxP8S37AYFku3hh4qiEif/4JFW5d+QKqdjTfBVQTRE34uOO3R07P6qmhemiePWWI
ERWa1cgf383MajvWFZZAkYc9Gq3SNoiCLJT3EWYRER/niYU2qnJOR8NsGJW5oPJx
PnmZyR3Tn86QN8tfn1/14mAx962bW9km4q6hz+9t9MYfz2/f4dyJjo3u6wAA3qeb
Zvn8HQrZjChqvQ/ryTd7yLxco/F7bUbtsjGC4hPlXNKdw6O3Gzy5HqmYtTa0Zc9I
5w1zNkoI7+ACQr3nhMKEL0EKwdHSdCreynOjsdr3BRTr2EK9Jeu1y80GDDQOec0z
B2ewl4C75fSrwLiG8/H3KsMFPcJh96J41G+JnMcrNIx8YqyMHksvVV6lAnlxC8hn
RzR4sgKkQ0A/rr5bPAIEQ5uOCiv5ZPTXGC89lat+acVi6koVGG01GqxwKTg3dOMy
lZzRMXjzdH4qJ3TNw5P+kRDU3nik+69Rx6nUnWBLPTkD77C5KU5q879iZShsdeSn
iST9/r0RAWWHut8xVRDSFJUk/dIHt+q0wyrs3yVrp0o1OpPo507FUmDH0jd41EtY
k3Dm1wo4SOyvoXloJTTrTc9aAcZREY4NfCKszo0v3t67uSf0RbTe8Vl1mJqkukhU
vyU/TI4STf2PnTrXboD3FOCyjU/3OOYfGFvTslr19Y8YoCBHBfBjo97/DruumToF
UmeaficW9Jeh/zub7F1GLHVaPcUeKUkxsOQPoMfcuC0BZijwzQePFTJoOVvLJD9x
Dk3pgjOr6ajSQ38Z+fm91dosntIf8FxYkcQrEojRxb3dAd5tPP5t8X0wuNu+KJmd
g7siGYBiOBmOh81tEQtf36BqEk6EZasWy5vJJTLvSARrKbqBU0+0Kf/Dv9Te7OL5
UIaY39SFRizOkpXID+lqEAGX2LwVQ7MrLQK1ycyfrVQ6aVW70ykMYxMVc0SKCqj/
ArX90N06+K/2xW5KTy0URgpnsLpX3dPtN+pW7S0TeudYhz6gdFJD9XeBq81j0TCy
fgycMTlutCL6MbV7+mwsv6T9Gm1RnirUBoq/CEYVql0xAmoIP27SUzaZMB5z+lQe
5sgiOjqONeu6Q3fsHN/iZa0L8sIps+0wsPFei9RlDP2ZHeFzASGbxNNaDy2i2d4V
ytKhjPm1T9ONb0w1NYoLMPUqR7K3jW9TlID0YCCyTWfX7Vhd9ME7MOq4cP7Euwl2
Z9h8wcCzfJd8hTDnB54l/uKrPb+MGiq+W6M0SoqNti6ShIJZuFfw72BbYxo/wgyD
3JKzgO0vC/eDf7Jpmm3eCN9PmlByWJRpEFw0DyLS8UhclEeiOko0W7830W38yt2e
DZVT+VkG4N8b8SsWlAzZIRhw+/ylAupuIyVvT+QOdo9meAjBECWR6bAu6lStsvux
Oox4l6cSBI1vmZqJp858QHDcLqFDt+ZTukisE8JRJoK7nKD9bxy1Os7vvf5CEdrT
eJQKiAMfd3OHSHCfALKq9nz3QBjZGemSFSHCHEwIYmKssxkVgP+6l01NGVQp0cMI
QbswMu74Is+3OPjogxoxndVTXlaQY/l1+8CBTyVzs/zmInxm2erYlUU19+38LUmi
murJx5bAsznv3ePTF4Ta2TFXsKozduK73dt6ebxnRMiqpBB5KXxHVBSLOaJZ2fHv
5UCypzJ38s+oBmczcYuKMLgcLjcdCdlccDTtkMIVcS+q6eaFKabMT0a4Q3B6TFqV
dmCePwzUYOb9XDgSc9ZpjdwiYkxVU0Yj1ChM6iTuv9OE2Vk6YxPDcnHvZ33fLWDG
ABz97nv1B0wzEQi5ZwO1dIrK/HvacvixwbuOlh0esw+2qhR5Affn8sKm9XrENJ5L
FqLtN8fJpf6X6RkzKC10Fs6/wr27a/PqhHOhm3N9EyZ9OXy5dTkLTOHU+wPKeBV6
0n1xzRxWLJcXEhzHfq40guAFk+3XW1CPNOLC2ObAQEDvFwyWX0l2z7wsKp9Gvquo
wC3hYNljjd260oFhcAR9ndD4D8V8lB7vTh1Q6gViiKM/iGqfCgUew2WRYYT8Gn2/
qoDXspokdFGsk3yoCfkIS38cN5uxr6jzO7JGLNsMl7eBuPyU9IjfDNLpb1UFrChd
TWqwydl5PsT6RWBqrS7Nf8lfXbOqUtZMJ/I5vPTwDs2blhuZk0LM7zaEPu+dL6m8
KcaVai0Lq+4ZwucHWP4w51S9NskcxvNo60uZmYbxDonJpmkStF+T/5xaw5oebqpB
qDAchuljScTgif5blXu3wv7I3lRcgivFzTgA8wue9IXi+vxqfYcjc75RbeMT/JtH
Itt77/kk5UUCCI4SUi0luP4hLCDk5/yASan7oX7rVGy7qOvZS/tdRl4ddhK3BExe
xui5HxE+laFL0dOBIH4MQxuzEQTQ7GiI07km7CWqLhl84TN5GKQOlRTBPFs4ADHK
w3IrO8g8LG1aQOdcbo4D2fNucUb16c5eO314D+wsfdWYCM11qaHhX/tCbcTcY+Ue
4H6Ug0xy4NJmw6OlMnq7rsSeJ7VtyacMxT1LG+Q/HERf4HaLXQtxCfJDVq8oU1M5
Izs7dT+OG0etWNBCV81yL9cv/3Uis9cq+mzfmLd7zdrKLnmcZ25SIBJ4ieWWe6/1
keTrMyR1QxLTrTWR+QIMrwvEfZRLnWD0ZmOgqLUbJNcSBkv7stzSCKDKLma3iHOS
KXvkAJ6Gc3rH9R1aVcCDHdFiHT6fbWHbpBeGE3UQ6ED4Q03E08IJvpF3l4uoXmc3
lWx8SNIlKfw2QtJMWOvPjyTevXB0CWb7+rTzWqweBRY97WVTWy8b8w4UUBOfDSIy
6ZmkZUH6IPQhKsm3Mo6I3HMHo7ms7nzx9J1lgJKPK4Ut9VBH2ykODcA5nIksPdk6
O+9Kbt8EJJNoH02goX1ipr0VzwPgdBFczHLDKS6wURzwtrKYXdQXzWfmHb92tl/B
ncLWBN4yvCZVIfuovo1XNQVipI2k9pL4oAlnGon8AyQ6e5UEDYrLtnhfU2p7sjbv
RwTJWH64fWO9VV67Zq6JU0kRt/IQnxguHXrZ0ADFgiSrxpn/XhDDZi3cuHggIe+v
5ksnf1ZVRMiYNUI3Y2KkTn6w4eg5XDzDuo6Vvqz0cQ+7w3SjiFEiJNNWy60Tl6rO
gRkSAWfyoxiKqSLttyvWgmAUuoJGWadGlIUE7uIZG3gC1s17kjtmns1tL6ejNaap
1St082obZGbDeL/T8i5018uEKtLdZ1pZq8U+lgIW5LAg+rvJ/QgyqglSXtmJj06d
gMsjpC+yPzfTXZz6ura/YIV4v4lYQ8K77WpIxzT9uBRHZOtl9mIqnBGASGZAB9Uo
JX0wyUvWDjuyGJWkkCu0XB3pfCgQi0spqPl/NNL+4hqZFuGeREmqZFVUTpUvA4Jb
ufN5E19sSvv1d0OdE+7RHQOaJ3ynB/mnoqk+8qQdiBJrWUC5UkdM9F4gPQpUyAKG
tkFA7OnAtWquxPHIIBLeoUP0oiZKw6Kf/4HXYHF1iGhsFRFa5dlNNO1AS7NGudMA
8gC+/n5wMr79i1hOII1slfrT+7NmPCs+4jTHjy3DtwOpp7w68dRyEISICu6Q5/qM
yS9elCoCapA+rp+7vosfUZgAosB8tmVbQPyXISwn0+fj0iiE1F4UBQ/yema1V1E+
uPQ4htNy5T5ByQVsQSRh0iUXYzeDjpwHiIRzrPlJOWCIUXcVUTJHRGI9jwIPZsU4
XjTQfkJa93B79/guFuRtiTfMKghq9OWqCXcSVEPnUt/61nnUxBR93yNrdqCcecZt
VAOsgJnKjkNwBbUE2KZfCJJOfc4t3RNqnpuUZkZptpbpw/xatUMhzHLwGx6hA27k
QE11tKJ966xWla+F2FzzlTGBj9dwbebnVQP3pTO4+Aek3Qi5CrPU8w3DDhYT/xh7
+Pck+DtuVdd+DtvadRdGxt/t6V09Rz/vK53yxx7XRafAgOH+os0a2j9+r1mDHDfa
WJLeYL84uNri3mpSionV90gcu2qrFvzFAPfPRvtCrtT+20uUay3Je7DqearU1wqy
7O+Ks2NfOBg/sSlQJA82U7v9/4fdlRPsqR9tkxSMbQm4ohYUgG0pS/HQ3P87V/mp
cYW9LXDHRgvR1EtxtJy/t+LC9HFrx2U+ZiuBV2MD5dyqhnGFONg4sii/wj/txjX+
l6buiqHkgfbHflBb6Gg+O+OhFqssaZ2j58D/huOzBVGvyzg1UAT31Paq498HSWEN
AgQGtGxhq1XPjX2oYEkBE8IhRw2g5ZW5jiwzMC2VP1rRXgzLfci/XQWwfrJ8NmzZ
LRRZXAOTqJSlLY6TCFQTfISY2b60gHPiHaZLnlPvsBHPTrT5Vlb+LQWo8Ni9vKFt
9tl96G1XiebxrxJpB8K52UgZsSfgn+Z8Bts/+SaZeF4NAWIj79VYXBZW0kgFOrfk
KTJsjQk8qGYCAZbCBBLQLrCFM5uABVbtekPUcI0eQR+okO9S8YMdOs4m7qng0Csh
NV8aVBA9BTuJTZQL+i92tYKGP3gxIme+aKxo/Rh//w6wy2LJ/48htixlMa5SYt/t
Fz2l3yPHj3s+b3uoMEFwo5P3xCh2WksKl/ftz/XuVtUO9EYHsgHnjZYNqLCp+yJk
tiENiUQ0Ky7yuGC4We8lePijrEyW9gji3XVFEAp2wdafR/JXKin7ir8NBQ984iDx
rTBL+BGpKAkebtaJ1Wp9yAIuagIjAiJ3BScvilPGfufHXRa2Nt4JevaalHDmTuu8
qlPuPxi2W9wzVcyYb+kYSTEoik1tkOsqkhhiUq6dJMAS1U2qNj/0V66mh+eHQKqg
1ATl4StO0D+v+C4W6u4TD3SMBNjWs2HYNohOID4Xc3OxFElUHHVIu7/NFCha65Py
wOw7zzU7ZGFEF0PuV83ajm3qAP+bYHSrkytC+FY06HCSn6ziio8YKkST+k1/C3rF
sTp4k1cyXwkn43s56IMhIjBZ1gldOfVmg5EGM8pXaZuQWT8ro48tlxFNxw+cIV71
QRWQ3WyDgdoSQJbZVx7Qe5Vgbc2Q44j9ESswsl3ZJjqM/aoqTDzjfgVSt+qi1RbT
+7WAVdICGPA7ABT4t3PkTzp2LBq8pII815neg7V5pKVzVJBP2Xwaru3QEzsUmAgb
GhP+VlKb0y/NDe0DGYLwbxYMmxvxYQtdUs6PznLDtLn9pHcvjeTDHl6e5WEQqz8E
+EHMI3U/1y4plv5xcyhPitQ+Dykdvh7d5vTd6bs+JnOyam6WNvHqVHaDmpesuhWb
SkNi5rp3UpHMyfP0oXKXmyqy6UAvINCDyMXhs5dQeTYcIu92gtrAajxw4s29wQV8
00yhb90rGc+G4NlAkxbszUDDTydnbnVs0Aw1OevNpL0oQt6jZBrEAid8NpNk2rwa
9/HfASdf0Q8i7O4kHe9BEEnSt+CaOpajU273TF6+q30s11e3FoIS9Ie/atJB/cuR
cCP//cbhZRSfMKn1kitYUlIoUkjb9sgKnGHX4w2f995Y0LQyV4PXUsiEtZDt/tcX
i8Umnwzc5RFyAgt0Aa7Af4CtyJtZCevyXj0P2/ZvAKq7kHMuAcx6w8WzaG8O4BDS
wCTqC0xF+vbp3jNMoPcvdPwhwguuAI3Fwxc0eW4KRS2QY4bpv46W007FZ1S5LSIs
gy9crusGHtP75eW1cX1Khjufw8dREXhREZyoUpB7dFFmdYJcb7p7pL1QaEIph9WZ
L29lYet1VrhP01P8B0Yf7zyieZw0p8xClZhNgW4e//81jBVXix/IrGv5/TKIsZDh
1LYSGOEGTWvkQkooJj4FgN9aQiYb1f/QdPTjra+B//lNxTbeuZXVCZIrpQjiUQUw
bZqF9214ZYmVQ8Pj8eQTMlNTQih5ueUCxsSBJ71Bvha7T8gl5ia0jrXHblu1E19S
lHf6gJfXZ60tudTKGb/WhLb6XvnH9V/bFyKeO/RoUku4whMFSpwHdiM/TUCXmBqW
GQfdj6LWLLSflRQP4W2RySUa65n04ouq6yv2wyMyETmo69UyKBgKnzE4B2njaIYz
RsasZZJtMKIc0M7qtlCDzCg9z/9sip631BKLce+1jACDN8xk40O7+P0DnZvidLZT
cQ3AjYVPin9OKLS5Y7I6oRXMMYeGMbWzYiBP+uO2GQg+AGsPE1RcABkDHVL8CiUR
5wtMXNoMkg4f6vJigVy7oI3iG8/xNvLGUucwL3z2IK76V8OQJEnOfDksyTZq2dgo
a23nHsfxGZ0au02TKZnh476G7uO1R2FWmp4SEyrizS2HJEVh1gL6yiXz6Jlh7eSL
EEHnHaGxAezAuZrpWzfG/hUGTL95VWgOFsc82SDbIdiO164xgSxj/FpEniczYU3G
JU5pTiyySS2f0E2yFzZkvIgrLN1Gfe710vsTXHKzxvIjfiBzkyFRBWmpS2euGLZE
pVzX7hlrTBtrGDvf4ct6dXv5R9P2PUptZojIosG5OwvM5vMwULQ3NaO/N8kfhtNb
ozyRMBnqAyOBnfnvL6GXYe5A1/B3U2kgVh+jTbyyeY1xTzYntIhNtO4e+1NHDSRO
M6deocHTk/2RRjXbLrrGQgHcad+keYQBRrxIOEzBn9Vn5dH5Ptgo55zZKGuLTRNf
E8JR4NO1TOyYt6X5nl884G+PUOaU+jZlV3AXZ/adkNMSSXp34E0jRUbNBncKtq/m
9vfSStSyHhmpoqDeWUXagmiG7ZQ6K3xLnIKxRY6m9n/4HVSXZ9Bmg+xXFz2XIi32
mhdyB6UFPJuDj0tQNjb/FYz2vJpiMvoYccixk2fhtOpRyxw/9qL9mHhB/gJSvdjY
GiV9uDlZJ7OtUsZIQjNi3f0gB8mnpXrsCqTDqS70cT9ToytcRgJ+W65T8h5QcR7z
I2GGnPa1k+I3LvOLAuCVBs9OXH135XYoBONzmmIdHCSiRL45XLBfOdcf9UrMG4a1
6x+OR3hG9duy1kw+Y8plFombnxUoG1vHB+/dISQl9TH3GDuhuPnEj/5psZIoWKBV
HRmhunecf8S9k4hj9+zv61Xpuaf6L712JXUF8gnMqeCIVMqUZSCOqT3sbc5dTrou
uDKh1LRG5p+1EFphwhHgaIOfSoUMseuxdtuZLuYvvjZkdSSsx6PWq+bfP6lNJYSt
V8bwyQyEDS22rzHXX54vB4fzlJXMyO5hQ/tOOq9PxJ5vZyuzbBfFlfdtFUyyVa3t
cijTAAk9/yweNarB2dVFpinXLpt6b8pwYJ+KQw2VaPNW9a3SNRVB1WtogwbAxUjs
16fkmZju78y7HnVI74aB1W05dBF2FLaQQ74BDN4/SFCq6qmDITb6+3AmChKmip2K
rF3WzmTE8LqVZ2PCntKhUbUBapRSH8g+4VKSJfaCIpv/tJBLEvgIOxkk7H0+Bk+y
LnaiKQBxaVljnoHuTmLGG3YvCPaMVVajOxEpVuvhNqcC6040qd90939I/dmkWESM
5fKWJg21fs+iQgyR1bIrg+q+l7W0GhBzFGrTzhzAKLcFml4RAbjlPVsZ0hXc3bIQ
t+jZIhoge/tkCDgT0/d2jjSa8/oso3KJ4oubjM5wTTxGAOO6TPHEHbRvv0z0ngBa
vIGd0vOMOVtnlRvyREw8TpLNqgTBRsqP5XT+yNDlFe4uweE9Dms/qtOBRwSzNZbw
kAUj9RH82pC8kNkVM7Aqaxx1+VE2ooTXnT9dENuHT0XBu8WRTNQrKZfMxmUh2L9o
Afjf6fEprIJ83cg9tJUp8prRGMt/7glWeY/R4YjqLmPc/i4mKs8kwiC6e233PZZ+
5iu2iowWCFmYpDHZvM/StYG6baOMtkDx53U83UunW5M/KYtHQHKPK5qBKwwN2vvq
n1V8l55+ywaHoNMCOmDNCALLHisa23KYupmwDroYUlI0vOEDWNGBr0K9WG677a25
a1LdNygdQITKVtDzJrX8rviqGn2LQskZ7mK4Bz7uH3mNGyK37KkZ3aSUps0n8tWm
HQhfjbTISMI2vfB7exObwtW4W0p22szoHjg9blms7eDMcZHozbU0gImvzDnxkf7T
6cphlMBCGE84bykxRq5Hl6Y8WRmx39KMkfq1gIowK2A5HpNZL9h/4i8UTCD7399/
UEcQDfgyv0wUc//oKp12tDxA9gkdDb6fR2JhNbpxnXsUnkrd8WKmxn0bXSxdYwOK
m73gyNSBQIoCwJxDDY4gwiOLpJAyoLU6/9ZrneRIe0nhH64eWg/cScj2veYMhRIV
RWrq+vGn/Btua07QGswMNHOGhE5yjaZndV7n0AcI4shtDjHUg+cvdSb6Ai2n1nGN
y0NG9vFJlZbx7MHkKU4f+VNCJZNSg+PMHkE0LMJasE1Z4pth3/lC2w1gS5GevvgY
W/QmkPmj5DsbcUiYMsoGmzEOBZbwD1hbih4bHujsDB0MAUhEQ8ChIMYg24m3XB9b
yo/PxGFJzJVBDALQh7xkCq7Q0j6QetjlKtou/go3oKRBWQLU0M1XIrceI9HHwjpS
luNUECk6+MzXSlclNsfCtZxj8iIC+H8KcqEeto0GJRP+RDJIfHkln0RIHnexzbSA
BARab5vRuK6xYBw0fjbdjb45RPh8SnIs9OAwaxtVKsMYUQUWBHdptriCr6uuSred
j3Vn1rSlWHhBR3bpe0Mihi+4ot6g3/Q/Dml/mhdOecnccQbAbdAErQZ2hLZsq6Of
9QsuayCeF6KTu9dZWWItyzvZ/lUHIu2Y4QpP+YLy7pGwfylWOGd0NMoOJBNVyeg+
mnIZeAQOJPvE8OheISX0QjC1fyfPmTqFIRKVNuD0ZsOY9xLMlK83bpLGqrpRmvK4
vFwFyLWBkuwy/NpyKzhvVtgwKx+G0cePMNeWfQ0mhUm1uNg97bfsuEPmCm6MbT3f
TVbBrl7iAIWlw111EgCQBxEiFCFXtgGDpi+59H9yhNmq4mZpM2PMsy3qI7koU3r6
SVzxP2VwIxLyPO9QGhAWpDbKw9qhw180U7r4ikHoUWkCOGvszFVqehrFmpLj8DR3
rCIYgQ1xSf0kSZIRPK/fHqRWW++huz7Il5vyV3yMyI0EIDkB6rpeO0VKoEUFwS4t
IIjA2p1ZWpKgmaw2ALWregkXq8vruu3C+KE6udyJcfH6O10+2uW4ZxeZstwrFXJv
CgLEHzoS3vTQoHL22aNoqjeRnx0H22POlJ8W1AoXk4Wn9MZE9beOGf1c+3o6ADS6
3tnuDJBdmWbGiueGMr35PFyIbwsajEUYpbZjn6QQ/GzxNTALuKHS6JKKywm2B94R
Ncrjrd12ORa4AmPKKHjrLFn6memejLbx0zdPJj3YGtGtxogNgjeeLVBQ5S9tzVic
Cbw80oDNTNB9RrUKj5wnqB2/MNeh4gsoshmcuvHYxKp2fmxxAOJ22ayILR+Kl904
xtAC3mDR4x99gkzFoJZ4qj9ZGGKZ8StS3CRDWQ8EgBWsN2udFP/3Fw5ZohvJXz9Y
P2q3F54nE6h27abmBBJbITRS7cl4+Ia78pAjRWd9PKSjeFzyOUtGUUWOHxJQox/2
sz/ib2Oz7cP7KxXYjoBuk5mhQgSCBDjPP6qJqvm+1il9rqyWD1q+KA4R5UIIF/u8
+vfgvUbXAxUbTq5uQaBphFA8OUf6vbJbnu3BZ1TQ28FnObnwvPRmsKMdUjR+YLgs
scmO05Xcz7WNJL5Oj4IAQXMYrrHeovF0YZYHLGloHEROd4+UKr8MVtmejvTbgwgX
NoBRzqxEKxdK7fVO5QnZMVoCay0T9Bas38zLxwk3B3LKz7LWsdC4gJfliNVi/nk7
+PGIapeZA1LaZ6XbZ+HP+zwlWqBZZwS7+vjHLjPJbqBb0L14MMUd1mMfEPTaxUYP
I5H8xkTqx9ni8RDzo7fCmsvbsJiCPAACyQRV7zki1CkW8zhr1+Yx8Jst+qS0Bcax
v+HoNX5rOYoRS5V8xqxWvXJAmvKNqyeIofx89vmwn11K4l6GBFFbkvr14qgwPbyF
EcBJq3qmW0JwKRcuoPdKmxeHDQ2nVsaw3pVPjQN4JfzWaNT5Yt8N9XQEy1VGw4DF
0J/OtZ5m8q+xRKrU1UFFU/Xa5tqnZMNL8m7CAz3Z6LHb3kUypYYYh0J1E5OKbw4c
AHBizHVNf31lhVY1YvmuB+BU9z3V20Ak3CyUV8oj6FOc0Wjt/U1nT5xQedgcmQUe
Tso3baTMY8+Nqw1UoFRMYuC2e0sdeFNG2twGhlhtHk7I3NgG4Y3QKaYuUHC8+OZ0
/Hle7itIc6Bud6vE8XQ2U+1c03Mt8cBiIzZnxPxOy77BfRh8VlGJ6r4H47lYZ7ui
JfydC/cGLDaS9d+h4QOSGsvSI4yodNOUZLra0ymI4AEj7s2vrc919VyMzBwXu1HB
qWmBDH9xED80uxi4bek0HydRCxUxsiMUs8hwQzYAjyJpRkm8cxecbYMiJCckH6Az
AhdFfp1C2FLfY36SGfWTprt3TkCHkLu9XvSdCFY1OeiV3R6Jl1AowpRKnCirMJ64
X3JYp5fqEVx6u8XzDr87t0Im4m/01WX8k46gK632Yr0tTD0tZlcdsZb3reEUaM8I
P8tlVZD0xScFY7ScgUK2DK5KYYmI/O00lAUtGSDmN5G8U7G/t9/F8Md/NMGRveBJ
VqkO3g8xMnM30sckHWwrWihiNhkoA4wHYhSlQfzCk2v/9F2HSDvrq9Ky/0pnd3xI
myimpDQOVSG0OYcci2ac4QEJTWSJeWPruEM4khjvToxjB1WKIxJ0m/GMiKesxIJu
K3eYOmeakt6+zzkTtrNDPpYbAMWU28zxp9sbhlWublspqpgPFVMlohDUJKtTecUQ
/G69uB1zOvUJ2XMrB0WQUvDVmrR3hgqdbZMNXIwKE2qiUhzEOnGzEBnmV9pObOAn
fXKewaMuEWikZanrBHJP1bKNNQNnQt0RWAtkgpcvUEtsYc/b6cPIEr8/JB64OPN1
iBLprgGTaSgqZxK9hBRAJvvshMLaPwnAeHwP5c0nOG2K8CxACrMXYoGTuUDImYSJ
+eo213ETz3jLF8ekazCsg9JQsRcEX0cYDCo/t/NGMECzBNbBZu1HVpJ7AFFxPe83
VoVlz1wXNN1Lhp2oh35+6g8fw6U2UhsSclTg2NZHlC/kimN2c+nHlgupE0zf65NQ
d8DrMVajG2CUa+lAinbPxR6hGx/0m8Y1qQGES1mKEcLqiFHacGIrDU+gWXTYPkyV
lmSqBKvbk9QdIyrreizSx6klRyUNT4aThXRKr9bzFzbWSI1ntl+Cz30AGGUsLcuo
VQu3V2mE9qWBpoh0EGX0281+2PznpIQgG+mNImKJbgGYezuo0qDIBWEJjZdszEqj
Zu94CarFaW/JC313I51N07lL7lpMlEjomhNgwuGX97vTD0I6YBp40fb7k4JUq92K
evxSurqgcpIYidpeY94egkGfADfLFEIm05ZGJ/VTR3OOWzpK9rfbPIF3ikCu/wrz
MgrlKKtFSPWxS0/CDYTQGVlw00ekx4i7En7KDD31N7CTdYXYPrg1vCA3BxD82LJ4
/7jUSutO0KeiwCxXorMowe68Tw70/7jfVSYmGLH5uAu9eMufrr2J6SjckJC/wWzj
R8vJM2CZhbHWpeo/a02ZFBrdJnUio1KkgJWMvCA+n7cyCJyru4LTtbXq/OQA5m2Z
BE/o97SUVh2P2DYZFXL/IdWkarvmWM2teWMtMNCpyl2lgcZ62zZMSp68ErsVvZbP
7vZkK7wW0vpn8IXX840IwTzasGdEc4IpCqySg7jAe3nkccx9678+EqLKUZVlaKBJ
ldyAQ4aFtD8LzTGjAttP6bSZ+CRomaD3A54X6tZD/+xCSgfosTDdovRhxvUtPVtp
6HJH/k21pgBgaxjp40Gr5alqHqGg/3d/yx9szKdZ6FiR+QgsPw6Q8XWOon+/2XiB
Ynt8ymSoe0OIePpPhyHuFS4sdNlzo264G7Nuu4B/iT4Vb1HRV10TrWxBDpDpBp7p
s2rharaG/byzcdW1N3UarM7mZ3t/oJnECl6UlXMnFU1wc6eHxm55shWZaRCWnxf3
lNGcCMZ10F4v5GiqEL85VIednx7JaRWcPaWCjjpFPLalyFaW3UgqUGzYG7SVWYv6
cHExhVnXsZEgTPKS4VGPbyfQSJ+yDaa7fDHiJNsj4BxjgMt97gSDubSuHnrZq9kJ
XW9Xy21S1aGvbg2THfg6BdWldsQ1i4OsSFBjNAtR+x3ci6Psk6KL3x1EZfK4efPK
UAnDoAosSoH4Zvk/LRE1bd6fCPwU3aoYDSXPSfLVQ9JXn6cPRXQXR93OJ7iaRinp
xk9c59551qJ/VIyPo5YILtjyqkYqqjoV1pZ23VfhAYAsTcMvO/aabP9mz9SH/9lG
p9zzlLAUhiT3uejEwlaBKQtSMP8HhMBYYfSYP8YNWHx7kW8aO4u2B3B/fUU/bf7k
dPi/sAczvVxninZer9UsEF1qSPVh7VP6NXpeCBR3NZptr4RQTSawzi7tnV7KVXO0
Nz+5geiX28kvqPiqc6SlJPS9hMi0od7EWM3m5Rz9bc3GisUqhOjVXwT8/aZRLegT
duBa0SWGcKNw6+rr7Rn7CK/pM0Une8thqKVvyHNa1kjDsX8vb2uvquMLkJ4fOxpJ
bCdtN/jyl62XexU2AvysmfnzQhbn1JWsUtcVs2hQb5WbR8+S+aRsiAmOUl6yGDjM
d/A6rPIGiV57CADaC++GQji1I4ntb8wIAvv4pXLYf/SzWSXt+rzX1aoxx+Ag138q
RI+XVSpWSjUaodRO1gjbYM5vQ0vWH3xl6fGCjNUO4yoMLY1hClG0vUqp/7KzGfN/
bNqB253gYm+Jy5SZ/p0/SgZUmysw+7wIpMuSDzsFKkAK2uUEY7PZ4LR+iQ8s/BNm
3d5xktUCfdYMqdC4X+HeeJywVgHu5foud0T/c67YgZYg4iHF38k8lHqG9cdOJ8w0
rIguqEFZNEqy6Ps73wwJzvN6DnJYiHvtNe4BA9TsN1JwtYjoNbeOqSwKc/ghEbIr
8A688j/UPIq4Jy0v3p0UiCcMTSKonyF9Ueb8s/DYWqB3niJO4AMWOgs9T+xszw3p
Z+KSQj89H2KQqylwYBwKgNSrt6+Ile4AeiQBqH74+wK4ow/VGnhPhI4859Sn5O/q
667Z5BOUuVgrraHjnmjf+4kzFJ2Vhiy4BbGiH3WzH3suzlb4e+n2GGwvXd2gYpoX
M1TPMr5uHMUDBeX6CHIsZT0P1F7sBm16xr+DbN6jYu8A2oSVPeykDNS+ByCTm5Oo
XkNfu/btabNayk+zqa8l7l5ADwj1S32y+DKyqtedc9kaMuEKeix+pTUFzqdxPfnh
yuIRNTHhx7yeYIdh95tb4PqJP1PeiALZTSTUjka9YUFxi5XWwfBZJHHujiXSdOMg
SF3uCNzcvfbLwY2T9m+Wo64wiz+3QUUIMk23npxT3yBYcEMP0DG0OAQSQVrxhh6c
BLG24UN0JjQGzGYLBSgc84aBfpabvMvBP0Aa8UxchSOKRtIlci+DoDKY2M8ZFe+B
asEC/2bEVNo1oEHbYo8frlf3gRO1qENuJN0SZ6cYRwzXIVGA+wTuumGyDzNjidcu
GibybJEqEZLOgoY3qXTdwt+V2T/HhRORWdjw5y8gJMBkmRyN/3+kJF4P7G3WnJAT
9WsqE6KeHutLGXRCXykb6Yv2crPSaAKzLPy6DSsy4l6tW7MsF2TXGBinIauun/HE
sxauRWMSu+m4UdMrQeIx2N7TivfdxQ00f0J7kHfQt6xi9IiOZEr1cJoLD6jjK7eU
B+MXiP5X66ym8cnrxD+8ERgUBlaH647XR9JbhU2cpetB8n/Hi5qoRlp8Rg4oPBlx
MAoKoxYFBHssIoJHAal92FlL+XSryFbja7mezpCmQiSv/6z8/y5H4yCa4KyHAxbf
YKgo/XfLhu0pWTYTgwNjpzxICgG3R50lP7fgnTr7+z5i3c6RTLOX7ft/ypko1LJy
JDwjiOVULKgJlee/wumLNKhJf7OcTzek6/GgsQY162D+FzOE0lOoyakFbThHMsbd
T+MF3iR9SQCQ0umoSIxOOgvI9WucH/CV0aLbdHGttCUNASYe/ucCVtxNbHEg8M6X
nfgmxmD3I5IwpAgkccLxsu17qPe9xuuIVy7mRRZT4kyZl61QjvI9WTec4qBfSZkN
JRskLV73jrbf7AARfRYJNumDMIb2z0qCK1S0jcvCqUA/xNWA1QOZH8FGXmJO0feO
U1LfhGcxX6CV3L+EqRJl6/iqhVeq8ldhgNEda99l0XPbjyfXKIDcFH0nJPCEe4zc
Py80FvVnUXyUcJdIAfk/dC6w8DxYC9l7LRScIm/FktU8yUsrf5gu3baw5Vnb4pNU
Mdsns7nDLsZZBJloPgChd2E8p/8J2T///cyyt4jcLLzEj8zxrWkx+wapM0GUhgw7
z/sXQMDgddJ6WTNGKfJ72u3FXh9wlL5KnXh18o4Nc87wcstvGYy0+apRJwEMVvz/
mk8+F3yuOt/PucDyUAMvkhpD2f5X34tDxtscs4bHVBY8GBQcSuSeloSV2jhB1/xI
E8crjNXT2zgF8H4VjBzWd1LXocAt6tuuAyX1XrR699/rtysLsv7E96xkYBfYP9li
+8umbCOED9xKHA7PAepBp7Cr+QIwFDqiDvMXJyvFi/+W57lBSUiXWZa3bMeMghIG
LDcEeOeZyAqD5xOscryQHrAqIZHy/lVyeCx1qEYCtusbIIWXdbNBWWN6IdRK52vz
iA3hK7UZWpLmg9Ml9NCNAEIjBTs1AcYyLH+0wLw/nAMOfg4WwUrGGLxXP/QZ78Zu
iLfVu0KtnDLri3MdmqCSlQHrOtDTf6kHTNlNZsGp6HA89EyJeFwrPERn+cTnefMG
c1gv1eEooh/7RRSgnMA3RaOrqGm8jHjYlTQxTvhC/Mzs812mQk8hWKa/cM0K6Ypl
U0uJ8F8wnH4YTl4j+HbkfUracdO7NFATPaAZezB1EBfju3sqzXKjHhHzM9Czx5v2
MzeiOlopyVrrj1fBf3vb37cJpiftXklYvxEOqnOdkZDwdlKUK7q9TX+/iHg4dJFA
YBLrRluckguv/ud3UFDF4pQZ8Hfw9yxAB+R7gD/aSvoBmoiRtysb1NGDxpXzF87o
wv4URv/mw5xnMh46ei2RfkGq7datUONJoj05j8oFr3JPNEl/L+dy+0jhFliFwjZX
IF0ElFtD/9XLgRhT50zNnNURnAXfyva0VjKTXbzkKxpXl7+cUkTU4K7M1704PGIW
vc17VmDdzxHX0kMTbbjJ4HL2QK1snPSpwPPW3pZkJEYjHIs5a2mYDBgEbcfEhZvJ
swVgsv1C5Eg6bxAFMzHDA+esWA5Qi/NWUU5zgLUsJ3W4YfyPQA0EYsIcd8tXdgHZ
l6nSZXKr3jp5ngVV0378n3oI54+HG9GclMuIVDY+PSnXJIIiGgNkp5VMMXqyWiW+
6FUmh7Jui7QmlbAKqp071aa+EgH6WfxQH4WkBweRvHzjb6uy/6xPEskfxZhyzIUU
wT4O31+159fD6Z9vNg/rMOBfn6YQo8w5Jmc/xZEO6CF9btloBLTueJoWTfRTXdMy
YIo6L6qgi57vojW3NRe7IPTs7RRHgEPop/ONzl7l2jbJD7j5xIwh4bjtn6mhI/PC
cTLnbMpoEa17He+HLjgIV8GZYB8CDfohUGB9kfph8HUINn3rWo6TQtMaYdx2vy1o
btRnoRTHkoITFr02rgZTliSUQX15Shhap9TR6ne9JmZpyP7mQv3s+AQu305dPQEq
UEOG8O6uX318YpYLMSRk2g1LMc5ustMfngEQRJeZ/00+g344df7frlu14Me7fBBU
McUQz/SjcWkkNGOzHT58Z8Sd3hZEbngIXQTTQ5GyKQSkXC85j40t/Tk8/Yr/S/xD
x93x/tk0QMQ4KWCIc0FoagH6RXOHn96sCJ7uBVrNy7A4kJrR0QlDbXc1lK93sLAd
iolpGBG7ks+vouCrSBgc/OSH+ZJ0rxiA+cIhaIBXEaVwGy6bGUJ/qWhjRMApa6hI
+yhnUbPs5Nxpw+vK0e+FuZncBxH064ogHi0pUfracToeHLsMPTMEAIlWGHN5NuzK
otig0li9ZRPcSqhOfFyQTrvZ18UWjwmDi/ik9DgD4Dmr5T//3czvVDrm3/XfCqkU
kV7JwXkEr4SAGoZJtFGSRyzoZnbMZfD2+EiU/2nA6FfcxhnzcQB7ejehNto8YEUC
wGfrrD1IpnnURSAtoXD0Rn0fSbi3bgmhzo/vikc3V0ySDVgsePyRXlk3+nMEbLjU
lZWRLbCUG26tKbJACfoDVuhu1n7aZZngAnObMJwMLeVtBsW916oCv8E1kcWHy1Vp
tjABSsVNJJI9f9xkB7vRXAYdxBuGuAnU9CbjNACSRNr/eoOjF42ErAb55Km+TCki
FRoFQZZ0hmjdY5356mrjEIz6oo/0ujtI8z5RTtZUSlqvuj7QmWKQs60na5nYhx2W
ndYJ9qBI4PAKrY6yZgA5dn3td5Fq41UxEAnHCu4Q7nRXo8E0PuXSpIlzGtwtaJqk
5jjqsUE/+OK8RRe1bCtNTyr2UQS0bZ6T+PYY+My3Nf7+v+zVvmnLGK9EDs65lnUF
N81oUbHLJGAB9un3+fDt7IyXfvWKDuAQDfkmJB/altuJ41nlOFwb1H9tQ8VBSTzA
XWge6FJGCDG2eIrWgwzERzN8ERDZzri4tfystk9LxTttW3EZucvh34BYXXXf57Nq
MP7Y40Jxpb2pT12p2C+KgZqKPTbEvJbzjoKo8NwoUFTmX1anjHEk7GOfjoa8MvDo
xEHpGuDyANdA6Hq0kz+JdRiZFGx+T1CrOfRvlXQVmlfoJQMWClV39mjRK4bj5LWv
91M4ZjAE57sqdjxkq0S8YgpxnqJr0hwRuTClR/0zzB1dUt05l7vkmIsxke4ZIwDn
1swcE7Ha6sAjusUe85UPwpmFtRvV5ZC/L6F38tyJv2ugC4SIXHV2NylH6jV3xyg3
fY9N/xrQ5zAKhi+Qdpgpljq5zy3mCKWnsQsQxwwW33UJejbxkUxTNVXR9e6pWjSm
sWJTb9N3mxkfwF/CzwyS54n2Xifr14KxXDscevIm3hytVdHNmpi+rhtZxU7fQ4ah
lGGOUCdBD+XH1KJRbOuyQqrRQuHAjcJA9NysUTHaa8HUuH0e35kUQRyF8PtrLkd3
32SKaC0t9LAl4PaTYFIPGx7Z8M4zsn24RqN2s5ZeRrfLyYcdFBqYm96c6mvsjFWS
qy1cSDHN5QKqJuf47MIOWA6e3v3M03wUFB0HYNGrKmpwxZ5CkFvBBJK3ZkHnKAF4
U0IRR+inWooDPIjmEcQWRVjX4io2eJQL5nrp7fzLU9v1iVwVRVGqNyqXGZlhU7bc
2jjteHYpYmch3zKP6SwkheET02O6wMQF0WyT4TUdV8RKhI6YmzGiZ9bL/vxcmU58
IQ7SS48AQ8VH4BNaUSS+HT5yqA8qCHZTsT/e6Fgu0BASzMAioJbPl8JxoE2oEy09
fGFvpglRvf08MQ+ICXulVoDUteJrPsfYshMYFdMBz6in2X5PsPuJrfofTgeBxG7w
nA3DYTjUqD+TbtZLQdlBx+x/kuC2JMMOldecgHN8dkcqmvDeVugy02ydQElsXR79
pWlXg1fxiQUei0+gtLMMb1fU67pWEyaWLQ9WK9BR/MOlYWQ8M+PDDZO0tjU4x0h9
INF8h3+6O2XdfbLOBObSn/SPx7NWl2etGDzjr+AJYpdUw0YnxraOtdvfXCmDkG7V
oTEBPSm/GnkLtomRn4IJyolvirrQtdLiD2ccSkNgKMEmlDR82m0e2oR/pZinbM/k
cCqLTHF9ln5IHjt2n9kuO3shUYMbNuC9tXvYyeeQRVuc5dNnHhxhGXnhVqDlecpF
8txxeImYXwebLAOxhWRC2RVDdjguo0Ie4t2CXp2eFoZoLnfBNrqbxQgwrYC9Per5
BIcFY/0coxRm2xcDLt98GK0cm95i1SKgxGyJoiRLNJEs5PJLdsmHTs4vycLuEwB1
+ovAwYBGpPTQD+/hokrwZg71BORqJdSTSu9A9mgvDETS4yQjyvuxu6N3UpPAyWmX
juuibzv/Rhe09xY8qI5zfLlDuwUtRWLQuF989FaP47bWZXUUa3jpdo7roc9XVeMN
NiiDWbORVw8U5aeYaClATFHTXUru/bq0XUVX/JlMkUDYvPlJWRahmX2+3hAWPNkP
m8dP/npKqgGjbOVtJ2j6lNqjrDAlg708H4iqjbbkZDiJ5GBWoEFuKSrcRU22si9k
L87IGokfBge+xOb8HJol3hr3Tp5uD7SWhSFcjy2UiqpUbwYEAfJpgfzVbdV9HG9P
CrGBnPW4AuDj/CNS+th8+SPtEqlcZbLoNB57/Ma0WHJGMBPaEeeWVCWaapUale37
3uloBd55M+2iufITENYzDJ/SkZtZGRHtkuvt46BtGsoCaxBCHmXkC8Ug9PoPacJI
/6WdToRA2lkfgos9ZGT26j3eGjRSw9UGL0G7v3TEiBoYmlmLu4RraSEXXkwAiUpe
VvMyUS9kfL9AqA9V3+xYlvEJVgxt9OfyRLmurVA3VPn/F+5HVhqdutTRg5z+bHVs
MU/O6z6deu+LtT+wh+b6fLMjO+ajQLsElqddhyPK3Y00fzGoPj7kbVXWpDGTyHMz
Gxc4kFMkgbLxTitV3rlXHF4d5xVaYCJCOjRDGT1YjhaGmilcdzJjxlWwOIgVak7J
i9VRY+rG6zO4GMqQpKhwqhYU1dKdx6CFjjRtYit53LewvrscAgGHzioK/E8aqQbr
uttiRuAEipMp9aVGBFSPhBGssqCcw+kzcLlJddYGcZDjlmVc8uTLIXcW5VMQAJ/k
1GTdafZqZ6SSQr2TNUJRWMLBtUonSRX5YMANO8+WX0ix7NuYgomQ56vgyxl+zBLp
fx19BxGLzGo3H0PQM8M2L6UwiSm2n870EwakQAE8YT0vELNcwYHHs+3gAtuUhZ4b
PWbKCZbGpPWesKoMx6Vc481u9fB6uuAXKKtQq/lpohHghyLVEf7runOHS30SbGNG
QYrXS8Rk/ZXUbMgz3VR+lg0wGsmF29+YiU5Sb6aA1+FlA3XEV9VjK4Z0MGlJ/PCl
rdVXZSOWF2UO+TAs6llji+OE8fY5TzzwiCrCkdtd3RHFh7LRBy8Eolm5pc19AZWL
VLGWI15AakitNXiW2yKNRKtmEz9rGggy/5cvAWuHNWRDKqNOq2TkO/flohLILEtx
D88r3pRNS5Zq+qNmhSqMKfaEZjfv20ogY5VBowTuDU7/5ti5PSZcLAmH7J5/+Ypd
Nc/AZ4XBzeVO3n9wH/lSgehWo792RUcmbXRY51NYnj43zA7YNoK4Da2VcJQsrU1g
RAcuh2Ypp6SZeWS6bF1e1bPNP895RGk/2h+nbEceRJPtPRddObK9b/GabEvDF0rs
jwfBpaoLRkmkNPazv6yfY8w+6aSN2dXFidWmS46PtD+lIlW7JKmE6FMSK5NufcxM
dfaVZoZgcxnd7EsvCXq5hwb77H9Fdd+9chSY8qLshFfAu3soO3/lmI3/11IxM0BG
kOTIU6t7DscsNtLMUE/a7Q4qMeZsnqbt+CafNBLm0Q+vB8bBEI3FGof26zA5nrD7
aZpMeKX2f9wAdrL8njQ3+PiTKf9LNOX/2PJYnHS925IF7An1YGnMgVykJkwGu+6Z
YcgsYt9qIrRrrgD6JUuYp6kKewDKusulvbjhmQk7RmoIHpYYx0ytyWh0IG0c09jy
FWt7odR8NKIMLCkgwjZkUYUlWTwBZMXDTQ7QyEw1XaCDax/Bq4sTi80m8JU1+FFZ
NYvGeR+MtIu5rLr7LKwXN0KLnPCy2TlyYdJMCktXcckIHlKnrbbjcBnXGc+pOZGd
oA1d7ZBLaDPVaiokYEm738syV1AG/q1+4fGiHJr81syL7c7sLkAcp+gys3u8APeV
kbWQN8TDJYSaMDY3KJubNuTdWWPdnvan5yS3If20D7uCikA5dPiMoL/6/B2CiOup
/O5YmgwlGDmIwQG6C70qRBCZ270ypgZuJkYdJZk6ySgjeQcS/Vb/VKpc2gECyrGK
H1OPp130S2edjUJzMDCkhjQpmDh1pJYIIIvsTc1vG+flxla1NjCLuLk8H1+sKT0J
lcmFekDIZHYM+L6w5n7OR1tiW55HtR+QSNRCTxWGTQ1wWziSuOYA9Fu8P28bKLz5
0Ak4m5Fnekwq1JrGBiK4znazolWOsZPQeCY7hnctXm+DcO0fUcTXZUEqfTaObLaM
PAn2CTIKzW9AraiHRve7HUb7TKVeeyEwJfHmkZvkFkUixQmNgX4Ae1zqosAnD6LG
S1//mj/28RQ0fS1r61rNJISWJETUJBSSgeAz/mIsPXOpAwdn8gizjI7g3reHvAsM
IrAmmP2JUY2Tb2pCNTZP5H+Uv4Jdr81l1IErS+GW7vn//nQ46sFNpkNk068gmQdP
eMQA7kRGPmnXohNosN8IeARdrsfuLYrxsYeAf5zfixJzUGW/KavVRYmKauOjapB1
JY8PtFhUxOCEk/PaeDHunRXxdxg7oST7R+iatIw9jsuiSmoZJxl08rK3et4DgE3w
sPHgQjpUDGyhogQ42acWsViwvqptJfTP+1CHbmXDdyipKtQeikveaNFZl8rMl2h3
t6Cq7wikQKu4eN1Jkhn1DdDf/q9fZDjcl1XGmt47ynYfiU6p62IcxgOrvSSlO5A5
Z8QUftMS8bXW0IPBMWDcDn4x+ovK5A5QWl2zdYNeh6moKELtKGAmlQomUAMDY5eQ
7Puhhr404dmjnggtWjJ0BLlF5BtzRbOs6cMOFZq1vz4J4etqcMSKIl7RhCerPX0J
3M4iRizwkc9jjr5goNrv0d5CWm2Pt+Q5WQhR7/Lp0qq/HenjaUaUVzcaIoJFnzXl
V5ruMvkxNjEWYizwX+N1QXrkwt94EDERNS7Drx/UyXQXznBfi+q2v5ycZ3LwSV/U
2QN44MHYsqjilX6NyiGzvSyqxgoAVRh+C+VXe8WuLBj+dlccDdKdNTQB/nGMgN0B
D8Q4w47wnb0mrQAaV8bFs7gPO3hydxwYCoqQBhTOFXqQY8IJSo9cElFb6YZzM+2F
DxInqM7iwFDkCYe0nNPk0xzJXt+dTANWmo5lJwRzEMMq1wbGB7XQyUKuiOAuECdI
3OYaMk4MlKAf6eAUzGW/oOml8ChZb1ajoQdtCA43lVvnVs6ow5Sc8FnnzZTjAzJS
e4Svx6kYYAIHCdIkwR/0yCmi3/SRGyqSuj+l1tiVcFsLsRzqVJZJjyQnuEa73rcS
zKQh7Bp57HceZ/0ivm+6wZlGCtYAxeUn7Jm6J1o5brrOIx7r3Vi9QtmETIe5LDi2
c+Jtvlw4uKBky9nMf6CrazkTDO4alR8zyodl9qhbkx83IsxRM+Cjpc9+eENQnDbf
of+XJBoCXj8vf00p9knJ3ZL1mm22QIGoxy7Ba4/j6ABDKqKTbVpijGkW9egKale0
6u5VsBFwmhMKKQumi3tA8UFFjnG7B+x3sz3alLU/dQ8En7SJXlQp67NS+Qk8S2AC
aGATgLEZq57VZ8MHyxp52pHeHd53kvRrSVq2DX4EfFGZeNQzQPKEu7rq8O+O9gnQ
MU/RU1YvNT2coqeV/PVtLmsUWPk+dhQvS7rL1GAp/RttSoEmvCZ5O4Lwsteodghu
Jq8eHUuns0QfPtSR3zyDxinu4ZhjEyOa+p/WkObdss0gdEQ/r/kgAav2irmOrAUC
KFFV7461xsGK94NaU2x1w5xzmfjlZjFpjNAcIBPnVa2kTkSooM5be0QCHPAkjB1D
lbCXpgWnf/lzYkcq4j6jJHNueYNktxEEFd9bg9xceAeuDyICVjRGm/6DqrywJ2nm
xwcSJI/OGLbpra0HPy9GF6GX/AuRIJWyHOijNvFcatRvB1mkdQ4bMv754XjNnbGW
tV5x5vgUdDvRC70HEwcwJvHCWVc1KN4/99hfOQtZTnmJvOTd91PmkMxN7KNR6qf9
QC+USeMph6LMrxDnJqSQ3vTRQJMsj1Ll6UbF+vgoKYs=
//pragma protect end_data_block
//pragma protect digest_block
JiOsrmr/aHun5dnMeA9kR1i+iWQ=
//pragma protect end_digest_block
//pragma protect end_protected
